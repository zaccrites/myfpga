
`ifndef MYFPGA_SVH
`define MYFPGA_SVH


`define NORTH   0
`define SOUTH   1
`define WEST    2
`define EAST    3

`define NORTHWEST   0
`define NORTHEAST   1
`define SOUTHWEST   2
`define SOUTHEAST   3


`endif


module slice (
    input logic i_ConfigDataIn,
    output logic o_ConfigDataOut,

);




shift_register8 config0 (

);

shift_register8 config1 (

);

shift_register8 config2 (

);



endmodule


module lut (

);

// Do something similar to Xilinx where they have a 6-input-1-output or 5-input-2-output?

mux8 mux(

);

endmodule


module logic_cell (

);

// two slices

endmodule
